interface top_interface_port;
logic clk;
logic rst_n;




endinterface