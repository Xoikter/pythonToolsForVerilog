interface test_interface_inner;




endinterface