class test_transaction extends uvm_sequence_item;



constraint con{


}
`uvm_object_utils_begin(test_transaction)


`uvm_object_utils_end
function new(string name = "test_transaction");
super.new();
endfunction
endclass
