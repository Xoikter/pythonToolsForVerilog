interface test_interface_port;
<<<<<<< HEAD
logic clk;
=======
>>>>>>> 51f05884d12d5605490827a74c95fc41601c853c
logic [3:0] a;
logic [3:0] b;
logic [4:0] c;




endinterface