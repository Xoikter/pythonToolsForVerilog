module topTB;
logic clk;
logic rst_n;
top topInst(
        .clk    (clk  ) ,//input   
        .rst_n  (rst_n));//input   
initial begin

end





endmodule
