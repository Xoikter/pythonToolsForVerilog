interface test_interface_port;
logic [3:0] a;
logic [3:0] b;
logic [4:0] c;
logic l;
logic as;




endinterface