module try(
	input clk,
	input rst_n,
	output reg q
);
reg p;

genvar i;
generate
	if (1) 
always@(posedge clk or negedge rst_n)

if (!rst_n) begin
q <= 0;
end
// else 
// q <= 0;
else
wire k = 1; 
endgenerate
endmodule