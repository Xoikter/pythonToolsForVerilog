interface top_interface_inner;




endinterface