interface test_interface;
test_interface_port ifo();
test_interface_inner ifi();




endinterface