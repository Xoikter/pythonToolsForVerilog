interface fifo_ctr_interface_inner;




endinterface