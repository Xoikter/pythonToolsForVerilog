interface top_interface;
top_interface_port if_o;
top_interface_inner if_i;




endinterface