interface test_interface;
<<<<<<< HEAD
test_interface_port ifo();
test_interface_inner ifi();


=======
// test_interface_port ifo();
// test_interface_inner ifi();
logic clk;
logic vld;
logic [3:0] a;
logic [3:0] b;
logic [4:0] c;
>>>>>>> 51f05884d12d5605490827a74c95fc41601c853c


endinterface