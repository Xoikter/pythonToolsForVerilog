interface test_interface;
// test_interface_port ifo();
// test_interface_inner ifi();
logic clk;
logic vld;
logic [3:0] a;
logic [3:0] b;
logic [4:0] c;


endinterface