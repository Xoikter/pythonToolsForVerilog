class top_transaction extends uvm_sequence_item;



constraint {


}
function new(string name = "top_transaction");
super.new();
endfunction
