class my_monitor extends uvm_monitor;

   virtual my_interface vif;
   uvm_active_passive_enum is_active = UVM_ACTIVE;
   uvm_analysis_port #(my_transaction)  ap;
   
   `uvm_component_utils(my_monitor)
   function new(string name = "my_monitor", uvm_component parent = null);
      super.new(name, parent);
   endfunction

   virtual function void build_phase(uvm_phase phase);
      int active;
      super.build_phase(phase);
      if(!uvm_config_db#(virtual my_interface)::get(this, "", "vif", vif))
         `uvm_fatal("my_monitor", "virtual interface must be set for vif!!!")
      ap = new("ap", this);      
      if(get_config_int("is_active", active)) is_active = uvm_active_passive_enum'(active);
   endfunction

   extern task main_phase(uvm_phase phase);
   extern task collect_one_pkt(my_transaction tr);
endclass

task my_monitor::main_phase(uvm_phase phase);
   my_transaction tr;
   //------------forever------//
   // while(1) begin
   //    tr = new("tr");
   //    collect_one_pkt(tr);
   //    ap.write(tr);
   // end

   //------------repeat-------//
   repeat(1) begin
      tr = new("tr");
      collect_one_pkt(tr);
      ap.write(tr);
   end


endtask

task my_monitor::collect_one_pkt(my_transaction tr);
      if(is_active == UVM_ACTIVE) begin

      end
      else begin

      end

endtask


