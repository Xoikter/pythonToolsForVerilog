interface top_interfac_port;
logic clk;
logic rst_n;




endinterface